`timescale 1ns / 1ps

/*
 * Copyright (c) 2023 Govardhan
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 */
module Data_Memory_tb;

   reg clk = 0; 
   reg WE;
   reg [31:0] A;
   reg [31:0] WD;
   wire [31:0] RD;

   always #5 clk = ~clk;

   Data_Memory Data_Memory_tb_inst (.clk(clk), .WE(WE), .A(A), .WD(WD), .RD(RD));

   initial begin
      WE = 0;
      A = 32'd10;
      WD = 32'd12345678;
      #10;
      WE = 1;
      #10;
      WE = 0;
      #10;
      A = 32'd20;
      WD = 32'd87654321;
      #10;
      WE = 1;
      #10;
      WE = 0;
      #10;
      $finish;
   end 

   initial begin
      $monitor("At time %d, RD = %h", $time, RD);
   end

endmodule
