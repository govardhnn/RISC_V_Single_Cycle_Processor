`timescale 1ns / 1ps
/*
 * Copyright (c) 2023 Govardhan
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 */
module PC_Mux_tb;

   reg [31:0] PC_Plus_4;
   reg [31:0] PC_Target;
   reg	      PCSrc;
   wire [31:0] PC_Next;

   PC_Mux PC_Mux_tb_inst (.PC_Plus_4(PC_Plus_4), .PC_Target(PC_Target), .PCSrc(PCSrc), .PC_Next(PC_Next));

   initial begin
      PC_Plus_4 = 32'd4;
      PC_Target = 32'd12345678;
      PCSrc = 0;
      #10;
      PCSrc = 1;
      #10;
      $finish;
   end 

   initial begin
      $monitor("At time %d, PC_Next = %d", $time, PC_Next);
   end

endmodule
